.title Amp

//Cascoded amp from [Sowlati 2002]

.include ../models/BFP620.lib
.include ../models/SMV2019079LF.lib
.include ../models/10pf0402.lib


Vsupply VCC 0 PULSE(0 4.0 20p 50p 10p 1ms 1ms)

Lsupply VCC D2 440NH

X1 D2 upper_base upper_E1 upper_E2 BFP620
X2 upper_E1 lower_base lower_E1 lower_E2 BFP620

C1 upper_base upper_base_ 0.1uF
Rb upper_base_ 0 50
Rb2 upper_base D2 1000

//X3 upper_base 0 10pf0402

Rgnd lower_E1 0 0

Lmatch D2 output_matched 2.2NH
Cmatch output_matched 0 0.4pF

Y1 output_matched 0 output 0 ymod
.MODEL ymod txl R=0.0236 L=0.306e-9 G=0.0001125 C=0.122e-12 length=10
//1.5 mm, 50-ohm trace on the 0.79mm substrates

Rout output 0 50

Lupper_bias upper_bias upper_base 50NH
Vupper_bias upper_bias 0 3

Rb3 lower_base lower_base_r 10
Vinp lower_base_r 0 SIN(0.7 0.7 8e9 0 0 0)

.control
//set num_threads=8

setcs DIOgradingCoeffMax=3.0
setcs DIOtDepCapMax = 2.0
tran 1p 300000ps uic
//uic?
plot D2 upper_E1
plot upper_base-upper_E1 lower_base
plot output
//plot collector
//plot b1 b2
//spec 0 15e9 3e7 v(collector)
//set specwindow = "blackman"
//plot mag(v(collector))
//set spectrum = mag(v(collector))

.endc

.end
