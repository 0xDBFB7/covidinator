.title Oscillator


.include ../models/BFP620.lib
.include ../models/SMV2019079LF.lib
.include ../models/10pf0402.lib


//Vsupply VCC 0 3.0
Vsupply VCC 0 PULSE(0 3.0 20p 5p 1p 1ms 1ms)

Lsupply VCC collector 440NH

X1 collector Base E1 E2 BFP620


//R1 collector in1 0 //0 ohm link
//R2 Base in2 0 //0 ohm link

//X2 collector in1 10pf0402
//X3 Base in2 10pf0402

Rbase_pulldown Base 0 10K //0 ohm link

R3 E1 0 0
R4 E2 0 0

P1 in1 in2 0 b1 b2 0 PLINE
.model PLINE CPL length={Len}
+R=1 0 1
+L={L11} {L12} {L22}
+G=0 0 0
+C={C11} {C12} {C22}
.param Len=6.5 Rs=0
.param Ceven_ground
.param Codd_
+ C11=0.3118p C12=-0.1797p C22=0.3118p
+ L11=0.3194NH L12=0.1887NH L22=0.3194NH

//length is in mm
//these are maxwellian matrix parameters.
//converted from physical parameters from wcalc
//coupled_microstrip.wc
//see Schutt‐Aine appnote,
//Relations Between Physical
//and Maxwellian Parameters
//(symmetric lines)

X4 b1 Varbias SMV2019079LF
X5 b2 Varbias SMV2019079LF
X6 0 Varbias SMV2019079LF
X7 0 Varbias SMV2019079LF
//C1 b1 0 0.31p
//C2 b2 0 0.31p

//varactors in series

R9 b1 0 10000
R8 b2 0 10000

R6 Varbias Vvaractor 20000
R7 Varbias Vvaractor 20000
Vcap Vvaractor 0 20.0

.ic v(Varbias) = 15


.control
//set num_threads=8
setcs DIOgradingCoeffMax=3.0
setcs DIOtDepCapMax = 2.0
tran 1p 100000ps uic
//uic?
//plot VCC Base
//plot collector
//plot b1 b2
//spec 0 15e9 3e7 v(collector)
//set specwindow = "blackman"
//plot mag(v(collector))
//set spectrum = mag(v(collector))

.endc

.end
