.title Amp

.include ../models/BFP620.lib
.include ../models/SMV2019079LF.lib
.include ../models/10pf0402.lib


Vsupply VCC 0 PULSE(0 5.0 20p 50p 10p 1ms 1ms)

Lsupply VCC D2 440NH

X1 D2 base E1 E2 BFP620

Re E1 0 25


Vbase base_bias 0 0.7

Rb base base_bias 50

Rbase base_ base 0
Cin input base_ 100pF

Vinp input 0 SIN(0 1 8e9 0 0 0)


Y1 D2 0 output 0 ymod
.MODEL ymod txl R=0.0236 L=0.306e-9 G=0.0001125 C=0.122e-12 length=10
//1.5 mm, 50-ohm trace on the 0.79mm substrates

Rout output 0 50

.control
//set num_threads=8

setcs DIOgradingCoeffMax=3.0
setcs DIOtDepCapMax = 2.0
tran 1p 300000ps uic
//uic?
plot D2 base
plot output
//plot collector
//plot b1 b2
//spec 0 15e9 3e7 v(collector)
//set specwindow = "blackman"
//plot mag(v(collector))
//set spectrum = mag(v(collector))

.endc

.end
