.title pore

Vsupply VCC 0 PULSE(0 1 20p 5p 1p 10ns 1us)


Rsolu VCC inp 100

Cmem1 inp m1 1NF
Rmem1 inp m1 10k

Rcore m1 m2 100

Rmem2 m2 0 10k
Cmem2 m2 0 1NF




.control
//set num_threads=8



setcs DIOgradingCoeffMax=3.0
setcs DIOtDepCapMax = 2.0
tran 1p 300000ps uic
//uic?
plot inp
plot (v(inp)-v(m1))
plot v(m2)

.endc

.end
