.title Oscillator


.include ../models/BFP620.lib
.include ../models/BFP540.lib
.include ../models/SMV2019079LF.lib
.include ../models/10pf0402.lib


Vsupply VCC 0 PULSE(0 2 20p 5p 1p 1ms 1ms)

Lsupply VCC collector 440NH

X1 collector Base E1 E2 BFP620

//LV1 Base Base_ 1.4NH
//X6 Base Base_ 10pf0402
X5 Base Base_ SMV2019079LF
X6 b___ Base_ SMV2019079LF
LV3 b___ 0 0NH
//C1 Base_ 0 0.3p


//LV2 collector collector__ 0.7NH
//X7 collector 0 10pf0402
//C2 collector__ 0 0.3p

X7 collector collector__ 10pf0402
X8 collector__ c__ SMV2019079LF
X9 c___ c__ SMV2019079LF
LV2 c___ 0 0NH
//X6 0 Base_ SMV2019079LF

Rbase_pulldown Base 0 10K //0 ohm link

Rc collector__ 0 10K //0 ohm link


Y1 collector 0 output 0 ymod
.MODEL ymod txl R=0.0236 L=0.306e-9 G=0.0001125 C=0.122e-12 length=5
//1.5 mm, 50-ohm trace on the 0.79mm substrates

Rout output 0 50

Y2 amp_C 0 amp_output 0 ymod
.MODEL ymod txl R=0.0236 L=0.306e-9 G=0.0001125 C=0.122e-12 length=5
Vamp_supply amp_supply 0 PULSE(0 5 50n 1n 1p 1ms 1ms)
Rsupply2 amp_supply amp_C 200
X2 amp_C amp_Base 0 0 BFP540ESD
Rbase1 amp_Base_ amp_Base 50
C2 output amp_Base_ 100pF
Rbase2 amp_Base amp_bias 150
Vbias amp_bias 0 0.6

Lem E1 E_ 440NH
Rem E_ E__ 1
Vem E__ 0 -1.0



Rem2 E1 E2 0


//X5 Base Varbias_2 SMV2019079LF
//X6 Varbias_2 0 10pf0402


R6 Base_ Vvaractor 10000
R7 collector__ Vvaractor 10000


.param varactor_bias_voltage = 15
Vcap Vvaractor 0 varactor_bias_voltage
//.ic v(Base_) = varactor_bias_voltage
//.ic v(Varbias_2) = varactor_bias_voltage


.control
//set num_threads=8



setcs DIOgradingCoeffMax=3.0
setcs DIOtDepCapMax = 2.0
tran 1p 300000ps uic
//uic?
plot output
plot amp_output
plot (v(amp_Base_)-v(amp_Base))/25
//plot collector
//plot b1 b2
//spec 0 15e9 3e7 v(collector)
//set specwindow = "blackman"
//plot mag(v(collector))
//set spectrum = mag(v(collector))

.endc

.end
